//-------------------------------------------------------------------------
//    Color_Mapper.sv                                                    --
//    Stephen Kempf                                                      --
//    3-1-06                                                             --
//                                                                       --
//    Modified by David Kesler  07-16-2008                               --
//    Translated by Joe Meng    07-07-2013                               --
//                                                                       --
//    Fall 2014 Distribution                                             --
//                                                                       --
//    For use with ECE 385 Lab 7                                         --
//    University of Illinois ECE Department                              --
//-------------------------------------------------------------------------


module  color_mapper ( input        [9:0] BallX, BallY, DrawX, DrawY, Ball_sizeX, Ball_sizeY, AlienX, AlienY,
                       output logic [7:0]  Red, Green, Blue );
    
    logic ship_on,alien_on;
	 
 /* Old Ball: Generated square box by checking if the current pixel is within a square of length
    2*Ball_Size, centered at (BallX, BallY).  Note that this requires unsigned comparisons.
	 
    if ((DrawX >= BallX - Ball_size) &&
       (DrawX <= BallX + Ball_size) &&
       (DrawY >= BallY - Ball_size) &&
       (DrawY <= BallY + Ball_size))

     New Ball: Generates (pixelated) circle by using the standard circle formula.  Note that while 
     this single line is quite powerful descriptively, it causes the synthesis tool to use up three
     of the 12 available multipliers on the chip!  Since the multiplicants are required to be signed,
	  we have to first cast them from logic to int (signed by default) before they are multiplied). */
	  
    int DistX, DistY, SizeX,SizeY;
	 assign DistX = DrawX - BallX;
    assign DistY = DrawY - BallY;
    assign SizeX = Ball_sizeX;
	 assign SizeY = Ball_sizeY;
	 
	 int DistX1, DistY1, SizeX1, SizeY1;
	 assign DistX1 = DrawX - AlienX;
    assign DistY1 = DrawY - AlienY;
    assign SizeX1 = Ball_sizeX;
	 assign SizeY1 = Ball_sizeY;
       
	  
    always_comb
    begin:Ship_on_proc
        //if ( ( DistX*DistX + DistY*DistY) <= (Size * Size) ) //ball
		  if(DistX>=0 && DistX<=SizeX &&DistY>=0&&DistY<=SizeY)  //square
            ship_on = 1'b1; 
        else 
            ship_on = 1'b0;
     end 
	  
	always_comb
	begin	:Alien_on_proc
	 //if ( ( DistX1*DistX1 + DistY1*DistY1) <= (Size1 * Size1) ) //ball
	 if(DistX1>=0 && DistX1<=SizeX1 &&DistY1>=0&&DistY1<=SizeY1) //square
            alien_on = 1'b1;
				else 
            alien_on = 1'b0;
	end
	
	always_comb
    begin:RGB_Display
        if ((ship_on == 1'b1)) 
        begin 
            Red = 8'hff;
            Green = 8'h55;
            Blue = 8'h00;
        end  
		  else if ((alien_on == 1'b1)) 
        begin 
            Red = 8'h00;
            Green = 8'h55;
            Blue = 8'h00;
        end 
        else 
        begin 
            Red = 8'h00; 
            Green = 8'h00;
            Blue = 8'h7f - DrawX[9:3];
        end      
    end 
    
endmodule
